module adder (a, b, s);
input [4:0] a,b;
output [4:0] s;
assign s = a + b;
endmodule
